module testb;halfadder_tb u1 (.co(co),.s(s),.a(a),.b(b)); halfadder u2 (.A(a),.B(b),.S(s),.CO(co)); endmodule